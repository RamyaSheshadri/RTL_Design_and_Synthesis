module mult2 (
    input [1:0] A,
    input [1:0] B,
    output [3:0] Y
);
    assign Y = A * B;
endmodule
